/* Dataflow style. */

module and_gate_dataflow (
    input a, b,
    output c
);
    assign c = a & b;
endmodule : and_gate_dataflow


/* End of file. */
