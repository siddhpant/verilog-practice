/* Dataflow style. */

module not_gate_dataflow (
    input a,
    output b
);
    assign b = ~a;
endmodule : not_gate_dataflow


/* End of file. */
